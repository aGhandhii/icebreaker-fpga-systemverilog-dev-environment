// Packages go in this directory
